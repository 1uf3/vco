* Created by KLayout

* cell TOP
.SUBCKT TOP
* net 15 Vout
* net 21 VDD
* net 27 GND
* cell instance $1 r0 *1 48.5,-18.9
X$1 27 5 20 19 18 17 21 21 21 21 21 26 25 24 10 23 11 9 8 1 3 1 11 9 8 3 12 1 9
+ 11 8 11 12 1 9 8 Inverter
* cell instance $2 r0 *1 334.2,10.5
X$2 1 Poly_cap
* cell instance $3 r0 *1 368.9,61.6
X$3 10 11 1 21 Pch
* cell instance $4 r0 *1 368.9,50.6
X$4 5 11 1 27 Nch
* cell instance $5 r0 *1 451.2,10.5
X$5 2 Poly_cap
* cell instance $6 r0 *1 485.9,61.6
X$6 14 3 2 21 Pch
* cell instance $7 r0 *1 485.9,50.6
X$7 7 3 2 27 Nch
* cell instance $8 r0 *1 446.9,61.6
X$8 13 2 12 21 Pch
* cell instance $9 r0 *1 446.9,50.6
X$9 6 2 12 27 Nch
* cell instance $12 r0 *1 260.7,-20.3
X$12 3 21 15 27 Buffer
* cell instance $13 r0 *1 490.2,10.5
X$13 3 Poly_cap
* cell instance $15 r0 *1 198.4,36.9
X$15 27 16 4 27 Nch$3
* cell instance $16 r0 *1 237.7,37.6
X$16 27 17 4 27 Nch$1
* cell instance $17 r0 *1 315.7,37.6
X$17 27 19 4 27 Nch$1
* cell instance $18 r0 *1 276.7,37.6
X$18 27 18 4 27 Nch$1
* cell instance $19 r0 *1 393.7,37.6
X$19 27 20 4 27 Nch$1
* cell instance $20 r0 *1 354.7,37.6
X$20 27 5 4 27 Nch$1
* cell instance $21 r0 *1 471.7,37.6
X$21 27 7 4 27 Nch$1
* cell instance $22 r0 *1 432.7,37.6
X$22 27 6 4 27 Nch$1
* cell instance $23 r0 *1 256.2,10.5
X$23 8 Poly_cap
* cell instance $24 r0 *1 295.2,10.5
X$24 9 Poly_cap
* cell instance $25 r0 *1 354.8,78.6
X$25 21 10 22 21 Pch$3
* cell instance $26 r0 *1 373.2,10.5
X$26 11 Poly_cap
* cell instance $27 r0 *1 412.2,10.5
X$27 12 Poly_cap
* cell instance $28 r0 *1 432.8,78.6
X$28 21 13 22 21 Pch$3
* cell instance $29 r0 *1 471.8,78.6
X$29 21 14 22 21 Pch$3
* cell instance $30 r0 *1 198.3,59.2
X$30 16 22 22 27 Nch$3
* cell instance $31 r0 *1 237.8,78.6
X$31 21 23 22 21 Pch$3
* cell instance $32 r180 *1 224.3,90.1
X$32 22 21 22 21 Pch$1
* cell instance $33 r0 *1 315.8,78.6
X$33 21 25 22 21 Pch$3
* cell instance $34 r0 *1 393.8,78.6
X$34 21 26 22 21 Pch$3
* cell instance $35 r0 *1 276.8,78.6
X$35 21 24 22 21 Pch$3
.ENDS TOP

* cell Poly_cap
* pin 
.SUBCKT Poly_cap 2
* device instance $1 r0 *1 14.8,10 CAP
C$1 2 1 1.12e-14 CAP
.ENDS Poly_cap

* cell Pch$3
* pin 
* pin 
* pin 
* pin 
.SUBCKT Pch$3 1 2 3 4
* device instance $1 r0 *1 4.5,4.5 PMOS
M$1 2 3 1 4 PMOS L=5U W=3U AS=6P AD=3P PS=10U PD=5U
* device instance $2 r0 *1 11.5,4.5 PMOS
M$2 1 3 2 4 PMOS L=5U W=3U AS=3P AD=3P PS=5U PD=5U
* device instance $3 r0 *1 18.5,4.5 PMOS
M$3 2 3 1 4 PMOS L=5U W=3U AS=3P AD=3P PS=5U PD=5U
* device instance $4 r0 *1 25.5,4.5 PMOS
M$4 1 3 2 4 PMOS L=5U W=3U AS=3P AD=6P PS=5U PD=10U
.ENDS Pch$3

* cell Nch$1
* pin 
* pin 
* pin 
* pin SUBSTRATE
.SUBCKT Nch$1 1 2 3 4
* net 4 SUBSTRATE
* device instance $1 r0 *1 4.5,4 NMOS
M$1 2 3 1 4 NMOS L=5U W=1U AS=4P AD=2P PS=8U PD=4U
* device instance $2 r0 *1 11.5,4 NMOS
M$2 1 3 2 4 NMOS L=5U W=1U AS=2P AD=2P PS=4U PD=4U
* device instance $3 r0 *1 18.5,4 NMOS
M$3 2 3 1 4 NMOS L=5U W=1U AS=2P AD=2P PS=4U PD=4U
* device instance $4 r0 *1 25.5,4 NMOS
M$4 1 3 2 4 NMOS L=5U W=1U AS=2P AD=4P PS=4U PD=8U
.ENDS Nch$1

* cell Buffer
* pin 
* pin 
* pin 
* pin SUBSTRATE
.SUBCKT Buffer 2 3 4 5
* net 5 SUBSTRATE
* cell instance $1 r0 *1 253.3,70.9
X$1 5 1 2 5 Nch
* cell instance $2 r0 *1 253.3,81.9
X$2 3 1 2 3 Pch
* cell instance $3 r0 *1 267.3,70.9
X$3 5 4 1 5 Nch
* cell instance $4 r0 *1 267.3,81.9
X$4 3 4 1 3 Pch
.ENDS Buffer

* cell Nch$3
* pin 
* pin 
* pin 
* pin SUBSTRATE
.SUBCKT Nch$3 1 2 3 4
* net 4 SUBSTRATE
* device instance $1 r0 *1 7,4 NMOS
M$1 2 3 1 4 NMOS L=10U W=2U AS=4P AD=2P PS=8U PD=4U
* device instance $2 r0 *1 19,4 NMOS
M$2 1 3 2 4 NMOS L=10U W=2U AS=2P AD=4P PS=4U PD=8U
.ENDS Nch$3

* cell Pch$1
* pin 
* pin 
* pin 
* pin 
.SUBCKT Pch$1 1 2 3 4
* device instance $1 r0 *1 7,6 PMOS
M$1 2 3 1 4 PMOS L=10U W=6U AS=12P AD=6P PS=16U PD=8U
* device instance $2 r0 *1 19,6 PMOS
M$2 1 3 2 4 PMOS L=10U W=6U AS=6P AD=12P PS=8U PD=16U
.ENDS Pch$1

* cell Inverter
* pin SUBSTRATE
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
.SUBCKT Inverter 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24
+ 25 26 27 28 29 30 31 32 33 34 35 36
* net 1 SUBSTRATE
* cell instance $1 r0 *1 203.4,69.5
X$1 6 36 26 1 Nch
* cell instance $2 r0 *1 242.4,69.5
X$2 5 35 25 1 Nch
* cell instance $3 r0 *1 281.4,69.5
X$3 4 34 24 1 Nch
* cell instance $4 r0 *1 359.4,69.5
X$4 3 33 23 1 Nch
* cell instance $5 r0 *1 320.4,69.5
X$5 2 32 22 1 Nch
* cell instance $6 r0 *1 359.4,80.5
X$6 12 27 17 7 Pch
* cell instance $7 r0 *1 281.4,80.5
X$7 13 28 18 8 Pch
* cell instance $8 r0 *1 242.4,80.5
X$8 14 29 19 9 Pch
* cell instance $9 r0 *1 320.4,80.5
X$9 15 30 20 10 Pch
* cell instance $10 r0 *1 203.4,80.5
X$10 16 31 21 11 Pch
.ENDS Inverter

* cell Pch
* pin 
* pin 
* pin 
* pin 
.SUBCKT Pch 1 2 3 4
* device instance $1 r0 *1 2.5,4.5 PMOS
M$1 2 3 1 4 PMOS L=1U W=3U AS=6P AD=6P PS=10U PD=10U
.ENDS Pch

* cell Nch
* pin 
* pin 
* pin 
* pin SUBSTRATE
.SUBCKT Nch 1 2 3 4
* net 4 SUBSTRATE
* device instance $1 r0 *1 2.5,4 NMOS
M$1 2 3 1 4 NMOS L=1U W=2U AS=4P AD=4P PS=8U PD=8U
.ENDS Nch
